module bcd7seg(
  input  [3:0] b,
  output reg [6:0] h
);

// 共阳极七段数码管段码定义:
//   a
//  ---
// f|   |b
//  ---  g
// e|   |c
//  ---  .dp
//   d

// 段码排列顺序: {g, f, e, d, c, b, a}  <-- 修改了这里
// 注意：0 表示点亮，1 表示熄灭 (因为是共阳极)

always @(*) begin
  case (b)
    4'b0000: h = 7'b1000000; // 0   <-- 修改了这里
    4'b0001: h = 7'b1111001; // 1
    4'b0010: h = 7'b0100100; // 2
    4'b0011: h = 7'b0110000; // 3
    4'b0100: h = 7'b0011001; // 4
    4'b0101: h = 7'b0010010; // 5
    4'b0110: h = 7'b0000010; // 6
    4'b0111: h = 7'b1111000; // 7
    4'b1000: h = 7'b0000000; // 8
    4'b1001: h = 7'b0010000; // 9
    4'b1010: h = 7'b0001000; // A
    4'b1011: h = 7'b0000110; // b
    4'b1100: h = 7'b1000110; // C
    4'b1101: h = 7'b0100001; // d
    4'b1110: h = 7'b0000111; // E
    4'b1111: h = 7'b0001110; // F
    default: h = 7'b1111111; // 默认情况，所有段熄灭
  endcase
end
endmodule